module nBit_Reg();
endmodule
