module multiplier();
endmodule
