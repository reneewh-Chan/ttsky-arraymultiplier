module fullAdder();
endmodule
