module nBit_register();
endmodule
